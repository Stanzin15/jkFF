class test;
    jk_env env_h;

    function new();
        env_h=new();
    endfunction 

    task run();
        env_h.run();
    endtask
endclass

